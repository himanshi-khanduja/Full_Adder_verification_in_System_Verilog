interface intf();
  
  logic a;
  logic b; 
  logic c;
  logic s;
  logic cout;
  
endinterface
